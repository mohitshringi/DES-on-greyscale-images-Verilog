`timescale 1ns / 1ns
module cbc_enc(final_cipher,input_grayscale_values,key,keyIV,clk);
output reg [1:8388608] final_cipher; 
input [1:64]  key;
input [1:64] keyIV;
input clk;                     
input [1:8388608] input_grayscale_values;

function [1:64] cypher(input [1:64] plain,input [1:64]  key);



   integer i;
   integer j;
   reg [1:7] IP[1:64];
   reg [1:7] PC1[1:56];
   reg [1:2] shift_left[1:16];
   reg [1:7] PC2[1:48];
   reg [1:64] new;
   reg [1:56] PC1perm;
   
   
   reg [1:32] L[0:16], R[0:16];
   reg [1:28] C[0:16], D[0:16];
   reg [1:56] cidi[1:16];
   reg [1:56] key1,key2,key3,key4,key5,key6,key7,key8,key9,key10,key11,key12,key13,key14,key15,key16;
   reg [1:48] K1,K2,K3,K4,K5,K6,K7,K8,K9,K10,K11,K12,K13,K14,K15,K16;
   reg [1:7] E[1:48];
   reg [1:48] T1;
   reg [1:4] S1[0:3][0:15];
   reg [1:4] S2[0:3][0:15];
   reg [1:4] S3[0:3][0:15];
   reg [1:4] S4[0:3][0:15];
   reg [1:4] S5[0:3][0:15];
   reg [1:4] S6[0:3][0:15];
   reg [1:4] S7[0:3][0:15];
   reg [1:4] S8[0:3][0:15];
   reg [1:6] P[1:32];
   reg [1:48] U1;
   reg [1:6] V11,V12,V13,V14,V15,V16,V17,V18;
   reg [1:2] Y11,Y12,Y13,Y14,Y15,Y16,Y17,Y18;
   reg [1:4] Z11,Z12,Z13,Z14,Z15,Z16,Z17,Z18;
   reg [1:4] W11,W12,W13,W14,W15,W16,W17,W18;
   reg [1:32] X1;
   reg [1:32] Q1;
   reg [1:64] result;
   reg [1:7] IP_inverse[1:64];
   

begin
IP[1] = 58;
			IP[2] = 50;
			IP[3] = 42;
			IP[4] = 34;
			IP[5] = 26;
			IP[6] = 18;
			IP[7] = 10;
			IP[8] = 2;
			IP[9] = 60;
			IP[10] = 52;
			IP[11] = 44;
			IP[12] = 36;
			IP[13] = 28;
			IP[14] = 20;
			IP[15] = 12;
			IP[16] = 4;
			IP[17] = 62;
			IP[18] = 54;
			IP[19] = 46;
			IP[20] = 38;
			IP[21] = 30;
			IP[22] = 22;
			IP[23] = 14;
			IP[24] = 6;
			IP[25] = 64;
			IP[26] = 56;
			IP[27] = 48;
			IP[28] = 40;
			IP[29] = 32;
			IP[30] = 24;
			IP[31] = 16;
			IP[32] = 8;
			IP[33] = 57;
			IP[34] = 49;
			IP[35] = 41;
			IP[36] = 33;
			IP[37] = 25;
			IP[38] = 17;
			IP[39] = 9;
			IP[40] = 1;
			IP[41] = 59;
			IP[42] = 51;
			IP[43] = 43;
			IP[44] = 35;
			IP[45] = 27;
			IP[46] = 19;
			IP[47] = 11;
			IP[48] = 3;
			IP[49] = 61;
			IP[50] = 53;
			IP[51] = 45;
			IP[52] = 37;
			IP[53] = 29;
			IP[54] = 21;
			IP[55] = 13;
			IP[56] = 5;
			IP[57] = 63;
			IP[58] = 55;
			IP[59] = 47;
			IP[60] = 39;
			IP[61] = 31;
			IP[62] = 23;
			IP[63] = 15;
			IP[64] = 7;
            
   for(i=1; i<=64; i=i+1)
   new[i]=plain[IP[i]];
   {L[0], R[0]} = new;
   
   PC1[1] = 57;
			PC1[2] = 49;
			PC1[3] = 41;
			PC1[4] = 33;
			PC1[5] = 25;
			PC1[6] = 17;
			PC1[7] = 9;
			PC1[8] = 1;
			PC1[9] = 58;
			PC1[10] = 50;
			PC1[11] = 42;
			PC1[12] = 34;
			PC1[13] = 26;
			PC1[14] = 18;
			PC1[15] = 10;
			PC1[16] = 2;
			PC1[17] = 59;
			PC1[18] = 51;
			PC1[19] = 43;
			PC1[20] = 35;
			PC1[21] = 27;
			PC1[22] = 19;
			PC1[23] = 11;
			PC1[24] = 3;
			PC1[25] = 60;
			PC1[26] = 52;
			PC1[27] = 44;
			PC1[28] = 36;
			PC1[29] = 63;
			PC1[30] = 55;
			PC1[31] = 47;
			PC1[32] = 39;
			PC1[33] = 31;
			PC1[34] = 23;
			PC1[35] = 15;
			PC1[36] = 7;
			PC1[37] = 62;
			PC1[38] = 54;
			PC1[39] = 46;
			PC1[40] = 38;
			PC1[41] = 30;
			PC1[42] = 22;
			PC1[43] = 14;
			PC1[44] = 6;
			PC1[45] = 61;
			PC1[46] = 53;
			PC1[47] = 45;
			PC1[48] = 37;
			PC1[49] = 29;
			PC1[50] = 21;
			PC1[51] = 13;
			PC1[52] = 5;
			PC1[53] = 28;
			PC1[54] = 20;
			PC1[55] = 12;
			PC1[56] = 4;
			
			for(i=1; i<=56; i=i+1)
        PC1perm[i] = key[PC1[i]];
        for(i=1; i<=28; i=i+1)
        C[0][i]=PC1perm[i];
        
        for(i=1; i<=28; i=i+1)
        D[0][i]=PC1perm[28+i];
        
        
        
   
      shift_left[1] = 1;
      shift_left[2] = 1;
      shift_left[3] = 2;
      shift_left[4] = 2;
      shift_left[5] = 2;
      shift_left[6] = 2;
      shift_left[7] = 2;
      shift_left[8] = 2;
      shift_left[9] = 1;
      shift_left[10] = 2;
      shift_left[11] = 2;
      shift_left[12] = 2;
      shift_left[13] = 2;
      shift_left[14] = 2;
      shift_left[15] = 2;
      shift_left[16] = 1;
      
      
      
      PC2[1] = 14;
			PC2[2] = 17;
			PC2[3] = 11;
			PC2[4] = 24;
			PC2[5] = 1;
			PC2[6] = 5;
			PC2[7] = 3;
			PC2[8] = 28;
			PC2[9] = 15;
			PC2[10] = 6;
			PC2[11] = 21;
			PC2[12] = 10;
			PC2[13] = 23;
			PC2[14] = 19;
			PC2[15] = 12;
			PC2[16] = 4;
			PC2[17] = 26;
			PC2[18] = 8;
			PC2[19] = 16;
			PC2[20] = 7;
			PC2[21] = 27;
			PC2[22] = 20;
			PC2[23] = 13;
			PC2[24] = 2;
			PC2[25] = 41;
			PC2[26] = 52;
			PC2[27] = 31;
			PC2[28] = 37;
			PC2[29] = 47;
			PC2[30] = 55;
			PC2[31] = 30;
			PC2[32] = 40;
			PC2[33] = 51;
			PC2[34] = 45;
			PC2[35] = 33;
			PC2[36] = 48;
			PC2[37] = 44;
			PC2[38] = 49;
			PC2[39] = 39;
			PC2[40] = 56;
			PC2[41] = 34;
			PC2[42] = 53;
			PC2[43] = 46;
			PC2[44] = 42;
			PC2[45] = 50;
			PC2[46] = 36;
			PC2[47] = 29;
			PC2[48] = 32;
      
        
        for(i=1; i<=16; i=i+1)
        begin
      if(shift_left[i]==2'b01)
      begin
      C[i][1]=C[i-1][28];
      for(j=1; j<=27; j=j+1)
      C[i][j+1]=C[i-1][j];
      D[i][1]=D[i-1][28];
      for(j=1; j<=27; j=j+1)
      D[i][j+1]=D[i-1][j];
      
       for(j=1; j<=28; j=j+1)
       cidi[i][j]=C[i][j];
       
       for(j=1; j<=28; j=j+1)
       cidi[i][j+28]=D[i][j];
       
      
      end  
      
      if(shift_left[i]==2'b10)
      begin
      C[i][1]=C[i-1][27];
      C[i][2]=C[i-1][28];
      for(j=1; j<=26; j=j+1)
      C[i][j+2]=C[i-1][j];
      D[i][1]=D[i-1][27];
      D[i][2]=D[i-1][28];
      for(j=1; j<=26; j=j+1)
      D[i][j+2]=D[i-1][j];
      
       for(j=1; j<=28; j=j+1)
       cidi[i][j]=C[i][j];
       
       for(j=1; j<=28; j=j+1)
       cidi[i][j+28]=D[i][j];
       
      
      
      end  
       
      
        end
        
        
        key1 = cidi[1];
        key2 = cidi[2];
        key3 = cidi[3];
        key4 = cidi[4];
        key5 = cidi[5];
        key6 = cidi[6];
        key7 = cidi[7];
        key8 = cidi[8];
        key9 = cidi[9];
        key10 = cidi[10];
        key11 = cidi[11];
        key12 = cidi[12];
        key13 = cidi[13];
        key14 = cidi[14];
        key15 = cidi[15];
        key16 = cidi[16];
        
        
        for(j=1; j<=48; j=j+1)
        K1[j]=key1[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K2[j]=key2[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K3[j]=key3[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K4[j]=key4[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K5[j]=key5[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K6[j]=key6[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K7[j]=key7[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K8[j]=key8[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K9[j]=key9[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K10[j]=key10[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K11[j]=key11[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K12[j]=key12[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K13[j]=key13[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K14[j]=key14[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K15[j]=key15[PC2[j]];
        
        for(j=1; j<=48; j=j+1)
        K16[j]=key16[PC2[j]];
      
      E[1] = 32;
			E[2] = 1;
			E[3] = 2;
			E[4] = 3;
			E[5] = 4;
			E[6] = 5;
			E[7] = 4;
			E[8] = 5;
			E[9] = 6;
			E[10] = 7;
			E[11] = 8;
			E[12] = 9;
			E[13] = 8;
			E[14] = 9;
			E[15] = 10;
			E[16] = 11;
			E[17] = 12;
			E[18] = 13;
			E[19] = 12;
			E[20] = 13;
			E[21] = 14;
			E[22] = 15;
			E[23] = 16;
			E[24] = 17;
			E[25] = 16;
			E[26] = 17;
			E[27] = 18;
			E[28] = 19;
			E[29] = 20;
			E[30] = 21;
			E[31] = 20;
			E[32] = 21;
			E[33] = 22;
			E[34] = 23;
			E[35] = 24;
			E[36] = 25;
			E[37] = 24;
			E[38] = 25;
			E[39] = 26;
			E[40] = 27;
			E[41] = 28;
			E[42] = 29;
			E[43] = 28;
			E[44] = 29;
			E[45] = 30;
			E[46] = 31;
			E[47] = 32;
			E[48] = 1;

S1[0][0] = 14;
			S1[0][1] = 4;
			S1[0][2] = 13;
			S1[0][3] = 1;
			S1[0][4] = 2;
			S1[0][5] = 15;
			S1[0][6] = 11;
			S1[0][7] = 8;
			S1[0][8] = 3;
			S1[0][9] = 10;
			S1[0][10] = 6;
			S1[0][11] = 12;
			S1[0][12] = 5;
			S1[0][13] = 9;
			S1[0][14] = 0;
			S1[0][15] = 7;
			S1[1][0] = 0;
			S1[1][1] = 15;
			S1[1][2] = 7;
			S1[1][3] = 4;
			S1[1][4] = 14;
			S1[1][5] = 2;
			S1[1][6] = 13;
			S1[1][7] = 1;
			S1[1][8] = 10;
			S1[1][9] = 6;
			S1[1][10] = 12;
			S1[1][11] = 11;
			S1[1][12] = 9;
			S1[1][13] = 5;
			S1[1][14] = 3;
			S1[1][15] = 8;
			S1[2][0] = 4;
			S1[2][1] = 1;
			S1[2][2] = 14;
			S1[2][3] = 8;
			S1[2][4] = 13;
			S1[2][5] = 6;
			S1[2][6] = 2;
			S1[2][7] = 11;
			S1[2][8] = 15;
			S1[2][9] = 12;
			S1[2][10] = 9;
			S1[2][11] = 7;
			S1[2][12] = 3;
			S1[2][13] = 10;
			S1[2][14] = 5;
			S1[2][15] = 0;
			S1[3][0] = 15;
			S1[3][1] = 12;
			S1[3][2] = 8;
			S1[3][3] = 2;
			S1[3][4] = 4;
			S1[3][5] = 9;
			S1[3][6] = 1;
			S1[3][7] = 7;
			S1[3][8] = 5;
			S1[3][9] = 11;
			S1[3][10] = 3;
			S1[3][11] = 14;
			S1[3][12] = 10;
			S1[3][13] = 0;
			S1[3][14] = 6;
			S1[3][15] = 13;
			S2[0][0] = 15;
			S2[0][1] = 1;
			S2[0][2] = 8;
			S2[0][3] = 14;
			S2[0][4] = 6;
			S2[0][5] = 11;
			S2[0][6] = 3;
			S2[0][7] = 4;
			S2[0][8] = 9;
			S2[0][9] = 7;
			S2[0][10] = 2;
			S2[0][11] = 13;
			S2[0][12] = 12;
			S2[0][13] = 0;
			S2[0][14] = 5;
			S2[0][15] = 10;
			S2[1][0] = 3;
			S2[1][1] = 13;
			S2[1][2] = 4;
			S2[1][3] = 7;
			S2[1][4] = 15;
			S2[1][5] = 2;
			S2[1][6] = 8;
			S2[1][7] = 14;
			S2[1][8] = 12;
			S2[1][9] = 0;
			S2[1][10] = 1;
			S2[1][11] = 10;
			S2[1][12] = 6;
			S2[1][13] = 9;
			S2[1][14] = 11;
			S2[1][15] = 5;
			S2[2][0] = 0;
			S2[2][1] = 14;
			S2[2][2] = 7;
			S2[2][3] = 11;
			S2[2][4] = 10;
			S2[2][5] = 4;
			S2[2][6] = 13;
			S2[2][7] = 1;
			S2[2][8] = 5;
			S2[2][9] = 8;
			S2[2][10] = 12;
			S2[2][11] = 6;
			S2[2][12] = 9;
			S2[2][13] = 3;
			S2[2][14] = 2;
			S2[2][15] = 15;
			S2[3][0] = 13;
			S2[3][1] = 8;
			S2[3][2] = 10;
			S2[3][3] = 1;
			S2[3][4] = 3;
			S2[3][5] = 15;
			S2[3][6] = 4;
			S2[3][7] = 2;
			S2[3][8] = 11;
			S2[3][9] = 6;
			S2[3][10] = 7;
			S2[3][11] = 12;
			S2[3][12] = 0;
			S2[3][13] = 5;
			S2[3][14] = 14;
			S2[3][15] = 9;
			S3[0][0] = 10;
			S3[0][1] = 0;
			S3[0][2] = 9;
			S3[0][3] = 14;
			S3[0][4] = 6;
			S3[0][5] = 3;
			S3[0][6] = 15;
			S3[0][7] = 5;
			S3[0][8] = 1;
			S3[0][9] = 13;
			S3[0][10] = 12;
			S3[0][11] = 7;
			S3[0][12] = 11;
			S3[0][13] = 4;
			S3[0][14] = 2;
			S3[0][15] = 8;
			S3[1][0] = 13;
			S3[1][1] = 7;
			S3[1][2] = 0;
			S3[1][3] = 9;
			S3[1][4] = 3;
			S3[1][5] = 4;
			S3[1][6] = 6;
			S3[1][7] = 10;
			S3[1][8] = 2;
			S3[1][9] = 8;
			S3[1][10] = 5;
			S3[1][11] = 14;
			S3[1][12] = 12;
			S3[1][13] = 11;
			S3[1][14] = 15;
			S3[1][15] = 1;
			S3[2][0] = 13;
			S3[2][1] = 6;
			S3[2][2] = 4;
			S3[2][3] = 9;
			S3[2][4] = 8;
			S3[2][5] = 15;
			S3[2][6] = 3;
			S3[2][7] = 0;
			S3[2][8] = 11;
			S3[2][9] = 1;
			S3[2][10] = 2;
			S3[2][11] = 12;
			S3[2][12] = 5;
			S3[2][13] = 10;
			S3[2][14] = 14;
			S3[2][15] = 7;
			S3[3][0] = 1;
			S3[3][1] = 10;
			S3[3][2] = 13;
			S3[3][3] = 0;
			S3[3][4] = 6;
			S3[3][5] = 9;
			S3[3][6] = 8;
			S3[3][7] = 7;
			S3[3][8] = 4;
			S3[3][9] = 15;
			S3[3][10] = 14;
			S3[3][11] = 3;
			S3[3][12] = 11;
			S3[3][13] = 5;
			S3[3][14] = 2;
			S3[3][15] = 12;
			S4[0][0] = 7;
			S4[0][1] = 13;
			S4[0][2] = 14;
			S4[0][3] = 3;
			S4[0][4] = 0;
			S4[0][5] = 6;
			S4[0][6] = 9;
			S4[0][7] = 10;
			S4[0][8] = 1;
			S4[0][9] = 2;
			S4[0][10] = 8;
			S4[0][11] = 5;
			S4[0][12] = 11;
			S4[0][13] = 12;
			S4[0][14] = 4;
			S4[0][15] = 15;
			S4[1][0] = 13;
			S4[1][1] = 8;
			S4[1][2] = 11;
			S4[1][3] = 5;
			S4[1][4] = 6;
			S4[1][5] = 15;
			S4[1][6] = 0;
			S4[1][7] = 3;
			S4[1][8] = 4;
			S4[1][9] = 7;
			S4[1][10] = 2;
			S4[1][11] = 12;
			S4[1][12] = 1;
			S4[1][13] = 10;
			S4[1][14] = 14;
			S4[1][15] = 9;
			S4[2][0] = 10;
			S4[2][1] = 6;
			S4[2][2] = 9;
			S4[2][3] = 0;
			S4[2][4] = 12;
			S4[2][5] = 11;
			S4[2][6] = 7;
			S4[2][7] = 13;
			S4[2][8] = 15;
			S4[2][9] = 1;
			S4[2][10] = 3;
			S4[2][11] = 14;
			S4[2][12] = 5;
			S4[2][13] = 2;
			S4[2][14] = 8;
			S4[2][15] = 4;
			S4[3][0] = 3;
			S4[3][1] = 15;
			S4[3][2] = 0;
			S4[3][3] = 6;
			S4[3][4] = 10;
			S4[3][5] = 1;
			S4[3][6] = 13;
			S4[3][7] = 8;
			S4[3][8] = 9;
			S4[3][9] = 4;
			S4[3][10] = 5;
			S4[3][11] = 11;
			S4[3][12] = 12;
			S4[3][13] = 7;
			S4[3][14] = 2;
			S4[3][15] = 14;
			S5[0][0] = 2;
			S5[0][1] = 12;
			S5[0][2] = 4;
			S5[0][3] = 1;
			S5[0][4] = 7;
			S5[0][5] = 10;
			S5[0][6] = 11;
			S5[0][7] = 6;
			S5[0][8] = 8;
			S5[0][9] = 5;
			S5[0][10] = 3;
			S5[0][11] = 15;
			S5[0][12] = 13;
			S5[0][13] = 0;
			S5[0][14] = 14;
			S5[0][15] = 9;
			S5[1][0] = 14;
			S5[1][1] = 11;
			S5[1][2] = 2;
			S5[1][3] = 12;
			S5[1][4] = 4;
			S5[1][5] = 7;
			S5[1][6] = 13;
			S5[1][7] = 1;
			S5[1][8] = 5;
			S5[1][9] = 0;
			S5[1][10] = 15;
			S5[1][11] = 10;
			S5[1][12] = 3;
			S5[1][13] = 9;
			S5[1][14] = 8;
			S5[1][15] = 6;
			S5[2][0] = 4;
			S5[2][1] = 2;
			S5[2][2] = 1;
			S5[2][3] = 11;
			S5[2][4] = 10;
			S5[2][5] = 13;
			S5[2][6] = 7;
			S5[2][7] = 8;
			S5[2][8] = 15;
			S5[2][9] = 9;
			S5[2][10] = 12;
			S5[2][11] = 5;
			S5[2][12] = 6;
			S5[2][13] = 3;
			S5[2][14] = 0;
			S5[2][15] = 14;
			S5[3][0] = 11;
			S5[3][1] = 8;
			S5[3][2] = 12;
			S5[3][3] = 7;
			S5[3][4] = 1;
			S5[3][5] = 14;
			S5[3][6] = 2;
			S5[3][7] = 13;
			S5[3][8] = 6;
			S5[3][9] = 15;
			S5[3][10] = 0;
			S5[3][11] = 9;
			S5[3][12] = 10;
			S5[3][13] = 4;
			S5[3][14] = 5;
			S5[3][15] = 3;
			S6[0][0] = 12;
			S6[0][1] = 1;
			S6[0][2] = 10;
			S6[0][3] = 15;
			S6[0][4] = 9;
			S6[0][5] = 2;
			S6[0][6] = 6;
			S6[0][7] = 8;
			S6[0][8] = 0;
			S6[0][9] = 13;
			S6[0][10] = 3;
			S6[0][11] = 4;
			S6[0][12] = 14;
			S6[0][13] = 7;
			S6[0][14] = 5;
			S6[0][15] = 11;
			S6[1][0] = 10;
			S6[1][1] = 15;
			S6[1][2] = 4;
			S6[1][3] = 2;
			S6[1][4] = 7;
			S6[1][5] = 12;
			S6[1][6] = 9;
			S6[1][7] = 5;
			S6[1][8] = 6;
			S6[1][9] = 1;
			S6[1][10] = 13;
			S6[1][11] = 14;
			S6[1][12] = 0;
			S6[1][13] = 11;
			S6[1][14] = 3;
			S6[1][15] = 8;
			S6[2][0] = 9;
			S6[2][1] = 14;
			S6[2][2] = 15;
			S6[2][3] = 5;
			S6[2][4] = 2;
			S6[2][5] = 8;
			S6[2][6] = 12;
			S6[2][7] = 3;
			S6[2][8] = 7;
			S6[2][9] = 0;
			S6[2][10] = 4;
			S6[2][11] = 10;
			S6[2][12] = 1;
			S6[2][13] = 13;
			S6[2][14] = 11;
			S6[2][15] = 6;
			S6[3][0] = 4;
			S6[3][1] = 3;
			S6[3][2] = 2;
			S6[3][3] = 12;
			S6[3][4] = 9;
			S6[3][5] = 5;
			S6[3][6] = 15;
			S6[3][7] = 10;
			S6[3][8] = 11;
			S6[3][9] = 14;
			S6[3][10] = 1;
			S6[3][11] = 7;
			S6[3][12] = 6;
			S6[3][13] = 0;
			S6[3][14] = 8;
			S6[3][15] = 13;
			S7[0][0] = 4;
			S7[0][1] = 11;
			S7[0][2] = 2;
			S7[0][3] = 14;
			S7[0][4] = 15;
			S7[0][5] = 0;
			S7[0][6] = 8;
			S7[0][7] = 13;
			S7[0][8] = 3;
			S7[0][9] = 12;
			S7[0][10] = 9;
			S7[0][11] = 7;
			S7[0][12] = 5;
			S7[0][13] = 10;
			S7[0][14] = 6;
			S7[0][15] = 1;
			S7[1][0] = 13;
			S7[1][1] = 0;
			S7[1][2] = 11;
			S7[1][3] = 7;
			S7[1][4] = 4;
			S7[1][5] = 9;
			S7[1][6] = 1;
			S7[1][7] = 10;
			S7[1][8] = 14;
			S7[1][9] = 3;
			S7[1][10] = 5;
			S7[1][11] = 12;
			S7[1][12] = 2;
			S7[1][13] = 15;
			S7[1][14] = 8;
			S7[1][15] = 6;
			S7[2][0] = 1;
			S7[2][1] = 4;
			S7[2][2] = 11;
			S7[2][3] = 13;
			S7[2][4] = 12;
			S7[2][5] = 3;
			S7[2][6] = 7;
			S7[2][7] = 14;
			S7[2][8] = 10;
			S7[2][9] = 15;
			S7[2][10] = 6;
			S7[2][11] = 8;
			S7[2][12] = 0;
			S7[2][13] = 5;
			S7[2][14] = 9;
			S7[2][15] = 2;
			S7[3][0] = 6;
			S7[3][1] = 11;
			S7[3][2] = 13;
			S7[3][3] = 8;
			S7[3][4] = 1;
			S7[3][5] = 4;
			S7[3][6] = 10;
			S7[3][7] = 7;
			S7[3][8] = 9;
			S7[3][9] = 5;
			S7[3][10] = 0;
			S7[3][11] = 15;
			S7[3][12] = 14;
			S7[3][13] = 2;
			S7[3][14] = 3;
			S7[3][15] = 12;
			S8[0][0] = 13;
			S8[0][1] = 2;
			S8[0][2] = 8;
			S8[0][3] = 4;
			S8[0][4] = 6;
			S8[0][5] = 15;
			S8[0][6] = 11;
			S8[0][7] = 1;
			S8[0][8] = 10;
			S8[0][9] = 9;
			S8[0][10] = 3;
			S8[0][11] = 14;
			S8[0][12] = 5;
			S8[0][13] = 0;
			S8[0][14] = 12;
			S8[0][15] = 7;
			S8[1][0] = 1;
			S8[1][1] = 15;
			S8[1][2] = 13;
			S8[1][3] = 8;
			S8[1][4] = 10;
			S8[1][5] = 3;
			S8[1][6] = 7;
			S8[1][7] = 4;
			S8[1][8] = 12;
			S8[1][9] = 5;
			S8[1][10] = 6;
			S8[1][11] = 11;
			S8[1][12] = 0;
			S8[1][13] = 14;
			S8[1][14] = 9;
			S8[1][15] = 2;
			S8[2][0] = 7;
			S8[2][1] = 11;
			S8[2][2] = 4;
			S8[2][3] = 1;
			S8[2][4] = 9;
			S8[2][5] = 12;
			S8[2][6] = 14;
			S8[2][7] = 2;
			S8[2][8] = 0;
			S8[2][9] = 6;
			S8[2][10] = 10;
			S8[2][11] = 13;
			S8[2][12] = 15;
			S8[2][13] = 3;
			S8[2][14] = 5;
			S8[2][15] = 8;
			S8[3][0] = 2;
			S8[3][1] = 1;
			S8[3][2] = 14;
			S8[3][3] = 7;
			S8[3][4] = 4;
			S8[3][5] = 10;
			S8[3][6] = 8;
			S8[3][7] = 13;
			S8[3][8] = 15;
			S8[3][9] = 12;
			S8[3][10] = 9;
			S8[3][11] = 0;
			S8[3][12] = 3;
			S8[3][13] = 5;
			S8[3][14] = 6;
			S8[3][15] = 11;







      for(i=1; i<=48; i=i+1)
        T1[i] = R[0][E[i]];
      
      U1 =K1^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      P[1] = 16;
			P[2] = 7;
			P[3] = 20;
			P[4] = 21;
			P[5] = 29;
			P[6] = 12;
			P[7] = 28;
			P[8] = 17;
			P[9] = 1;
			P[10] = 15;
			P[11] = 23;
			P[12] = 26;
			P[13] = 5;
			P[14] = 18;
			P[15] = 31;
			P[16] = 10;
			P[17] = 2;
			P[18] = 8;
			P[19] = 24;
			P[20] = 14;
			P[21] = 32;
			P[22] = 27;
			P[23] = 3;
			P[24] = 9;
			P[25] = 19;
			P[26] = 13;
			P[27] = 30;
			P[28] = 6;
			P[29] = 22;
			P[30] = 11;
			P[31] = 4;
			P[32] = 25;
     
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[1]=R[0];
      R[1]=L[0] ^ Q1;
      
      
      
       for(i=1; i<=48; i=i+1)
        T1[i] = R[1][E[i]];
      
      U1 =K2^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[2]=R[1];
      R[2]=L[1] ^ Q1;
      
      
      
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[2][E[i]];
      
      U1 =K3^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[3]=R[2];
      R[3]=L[2] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[3][E[i]];
      
      U1 =K4^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[4]=R[3];
      R[4]=L[3] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[4][E[i]];
      
      U1 =K5^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[5]=R[4];
      R[5]=L[4] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[5][E[i]];
      
      U1 =K6^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[6]=R[5];
      R[6]=L[5] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[6][E[i]];
      
      U1 =K7^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[7]=R[6];
      R[7]=L[6] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[7][E[i]];
      
      U1 =K8^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[8]=R[7];
      R[8]=L[7] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[8][E[i]];
      
      U1 =K9^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[9]=R[8];
      R[9]=L[8] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[9][E[i]];
      
      U1 =K10^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[10]=R[9];
      R[10]=L[9] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[10][E[i]];
      
      U1 =K11^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[11]=R[10];
      R[11]=L[10] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[11][E[i]];
      
      U1 =K12^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[12]=R[11];
      R[12]=L[11] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[12][E[i]];
      
      U1 =K13^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[13]=R[12];
      R[13]=L[12] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[13][E[i]];
      
      U1 =K14^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[14]=R[13];
      R[14]=L[13] ^ Q1;
      
      
      for(i=1; i<=48; i=i+1)
        T1[i] = R[14][E[i]];
      
      U1 =K15^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[15]=R[14];
      R[15]=L[14] ^ Q1;
      
      
      
       for(i=1; i<=48; i=i+1)
        T1[i] = R[15][E[i]];
      
      U1 =K16^T1;
      
      for(i=1; i<=6; i=i+1)
        V11[i] = U1[i];
        for(i=7; i<=12; i=i+1)
        V12[i-6] = U1[i];
        for(i=13; i<=18; i=i+1)
        V13[i-12] = U1[i];
        for(i=19; i<=24; i=i+1)
        V14[i-18] = U1[i];
        for(i=25; i<=30; i=i+1)
        V15[i-24] = U1[i];
        for(i=31; i<=36; i=i+1)
        V16[i-30] = U1[i];
        for(i=37; i<=42; i=i+1)
        V17[i-36] = U1[i];
        for(i=43; i<=48; i=i+1)
        V18[i-42] = U1[i];
        
      Y11[1]=V11[1];
      Y11[2]=V11[6];
      Z11[1]=V11[2];
      Z11[2]=V11[3];
      Z11[3]=V11[4];
      Z11[4]=V11[5];
      
       Y12[1]=V12[1];
      Y12[2]=V12[6];
      Z12[1]=V12[2];
      Z12[2]=V12[3];
      Z12[3]=V11[4];
      Z12[4]=V12[5];
      
       Y13[1]=V13[1];
      Y13[2]=V13[6];
      Z13[1]=V13[2];
      Z13[2]=V13[3];
      Z13[3]=V13[4];
      Z13[4]=V13[5];
      
       Y14[1]=V14[1];
      Y14[2]=V14[6];
      Z14[1]=V14[2];
      Z14[2]=V14[3];
      Z14[3]=V14[4];
      Z14[4]=V14[5];
      
       
      
       Y15[1]=V15[1];
      Y15[2]=V15[6];
      Z15[1]=V15[2];
      Z15[2]=V15[3];
      Z15[3]=V15[4];
      Z15[4]=V15[5];
      
       Y16[1]=V16[1];
      Y16[2]=V16[6];
      Z16[1]=V16[2];
      Z16[2]=V16[3];
      Z16[3]=V16[4];
      Z16[4]=V16[5];
      
       Y17[1]=V17[1];
      Y17[2]=V17[6];
      Z17[1]=V17[2];
      Z17[2]=V17[3];
      Z17[3]=V17[4];
      Z17[4]=V17[5];
      
      Y18[1]=V18[1];
      Y18[2]=V18[6];
      Z18[1]=V18[2];
      Z18[2]=V18[3];
      Z18[3]=V18[4];
      Z18[4]=V18[5];
      
      W11=S1[Y11][Z11];
       W12=S2[Y12][Z12];
        W13=S3[Y13][Z13];
         W14=S4[Y14][Z14];
          W15=S5[Y15][Z15];
         W16=S6[Y16][Z16];
          W17=S7[Y17][Z17];
           W18=S8[Y18][Z18];
           
      for(i=1;i<=4;i=i+1)
      X1[i]=W11[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+4]=W12[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+8]=W13[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+12]=W14[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+16]=W15[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+20]=W16[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+24]=W17[i];
      
      for(i=1;i<=4;i=i+1)
      X1[i+28]=W18[i];
      
      
      
     for(i=1;i<=32;i=i+1)
     Q1[i]=X1[P[i]];
      
        
      L[16]=R[15];
      R[16]=L[15] ^ Q1;
      
      
      
       //cipher=R[16];
    
    
    
    for(i=1;i<=32;i=i+1)
    result[i]=R[16][i];
    
    for(i=1;i<=32;i=i+1)
    result[i+32]=L[16][i];
    
   
   
   
   IP_inverse[1] = 40;
			IP_inverse[2] = 8;
			IP_inverse[3] = 48;
			IP_inverse[4] = 16;
			IP_inverse[5] = 56;
			IP_inverse[6] = 24;
			IP_inverse[7] = 64;
			IP_inverse[8] = 32;
			IP_inverse[9] = 39;
			IP_inverse[10] = 7;
			IP_inverse[11] = 47;
			IP_inverse[12] = 15;
			IP_inverse[13] = 55;
			IP_inverse[14] = 23;
			IP_inverse[15] = 63;
			IP_inverse[16] = 31;
			IP_inverse[17] = 38;
			IP_inverse[18] = 6;
			IP_inverse[19] = 46;
			IP_inverse[20] = 14;
			IP_inverse[21] = 54;
			IP_inverse[22] = 22;
			IP_inverse[23] = 62;
			IP_inverse[24] = 30;
			IP_inverse[25] = 37;
			IP_inverse[26] = 5;
			IP_inverse[27] = 45;
			IP_inverse[28] = 13;
			IP_inverse[29] = 53;
			IP_inverse[30] = 21;
			IP_inverse[31] = 61;
			IP_inverse[32] = 29;
			IP_inverse[33] = 36;
			IP_inverse[34] = 4;
			IP_inverse[35] = 44;
			IP_inverse[36] = 12;
			IP_inverse[37] = 52;
			IP_inverse[38] = 20;
			IP_inverse[39] = 60;
			IP_inverse[40] = 28;
			IP_inverse[41] = 35;
			IP_inverse[42] = 3;
			IP_inverse[43] = 43;
			IP_inverse[44] = 11;
			IP_inverse[45] = 51;
			IP_inverse[46] = 19;
			IP_inverse[47] = 59;
			IP_inverse[48] = 27;
			IP_inverse[49] = 34;
			IP_inverse[50] = 2;
			IP_inverse[51] = 42;
			IP_inverse[52] = 10;
			IP_inverse[53] = 50;
			IP_inverse[54] = 18;
			IP_inverse[55] = 58;
			IP_inverse[56] = 26;
			IP_inverse[57] = 33;
			IP_inverse[58] = 1;
			IP_inverse[59] = 41;
			IP_inverse[60] = 9;
			IP_inverse[61] = 49;
			IP_inverse[62] = 17;
			IP_inverse[63] = 57;
			IP_inverse[64] = 25;

			for(i=1; i<=64; i=i+1)
       cypher[i]=result[IP_inverse[i]];
       
end
endfunction

 reg [1:64] temp_plain;  
 reg [1:64] first;
  
 integer k=1;
  integer l=1;
  
  /*
    ******
    ******
    CHANGE FILE LOCATION IN THE VARIABLE BELOW AS PER YOUR PC
    ******
    ******
    */ 
  integer output_file;
  initial output_file=$fopen("D:/I-CHIP_2bits/cbc_enc_out.txt");
  
  always @ (posedge clk, negedge clk)                        
  begin                                        
   temp_plain=input_grayscale_values[k+:64];  
    if(k==1)
    begin
     first = temp_plain^keyIV;
     final_cipher[1:64]=cypher(first,key);
     
    $fwrite(output_file,"%b",final_cipher[1:64]);
     k=k+64;
     end      
   
    else 
    begin
    if(k>=8388608) begin $fclose(output_file);
    $finish;
    end
     first = temp_plain ^ final_cipher[l+:64];  
     final_cipher[k+:64]=cypher(first,key); 
     
    $fwrite(output_file,"%b",final_cipher[k+:64]);
    
     k=k+64;l=l+64;
    end     
    
  end 
  
endmodule
